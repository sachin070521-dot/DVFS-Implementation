`timescale 1ns / 1ps
module dfs_alu_top (
    input  wire        clk_100mhz,   // 100 MHz Basys-3 clock
    input  wire        rst,

    // ALU control (can come from switches / testbench)
    input  wire        alu_en,
    input  wire [2:0]  alu_op,
    input  wire [31:0] alu_a,
    input  wire [31:0] alu_b,

    // Debug output
    output wire led0,   // blink (frequency effect)
    output wire led1,   // dfs_sel[0]
    output wire led2,
    output wire led3   // dfs_sel[1]
  );
    // =====================================================
    // 1. Clock Divider
    // =====================================================
    wire clk_div2, clk_div4, clk_div8;

    clock_divider u_div (
        .clk_in   (clk_100mhz),
        .rst      (rst),
        .clk_div2 (clk_div2),
        .clk_div4 (clk_div4),
        .clk_div8 (clk_div8)
  
   );
    // =====================================================
    // 2. DFS Clock Select (AUTOMATIC)
    // =====================================================
    wire [1:0] dfs_sel;
    wire       dfs_clk;

    assign dfs_clk =
        (dfs_sel == 2'b10) ? clk_div2  :   // HIGH activity  -> f/2
        (dfs_sel == 2'b01) ? clk_div4  :   // MED activity   -> f/4
                             clk_div8 ;   // LOW activity   -> f/8

    // =====================================================
    // 3. ALU
    // =====================================================
    wire [31:0] alu_y;
    wire        alu_valid;

    alu_32bit u_alu (
        .clk   (dfs_clk),
        .rst   (rst),
        .en    (alu_en),
        .op    (alu_op),
        .a     (32'd4500),
        .b     (32'd200),
        .y     (alu_y),
        .valid (alu_valid)
    );

    // =====================================================
    // 4. Activity Monitor
    // =====================================================
    wire [15:0] activity;

    activity_monitor u_activity (
        .clk       (dfs_clk),
        .rst       (rst),
        .alu_valid (alu_valid),
        .activity  (activity)
    );

    // =====================================================
    // 5. DFS Controller
    // =====================================================
    dfs_controller u_dfs_ctrl (
        .clk      (clk_100mhz),   // control logic runs on base clock
        .rst      (rst),
        .activity (activity),
        .dfs_sel  (dfs_sel)
    );

    // =====================================================
    // 6. LED Debug (Human-visible DFS effect)
    // =====================================================
    reg [25:0] led_cnt;
    reg        led_blink;

    always @(posedge dfs_clk or posedge rst) begin
        if (rst) begin
            led_cnt   <= 0;
            led_blink <= 0;
        end else begin
            led_cnt <= led_cnt + 1;
            if (led_cnt == 26'd0)
                led_blink <= ~led_blink;
        end
    end

    assign led0 = led_blink;              // Blink = DFS clock speed
assign led1 = dfs_sel[0] & led_blink; // MED indicator
assign led2 = dfs_sel[1] & led_blink; // HIGH indicator
assign led3 = 1'b0; 
assign led4 = (activity[15:14] != 2'b00);   // very low → low
assign led5 = (activity[15:13] != 3'b000);  // low → medium
assign led6 = (activity[15:12] != 4'b0000); // medium → high
assign led7 = (activity[15:11] != 5'b00000);// very high                  // unused
endmodule
